//////////////////
// Memory stage //
//////////////////

module kamacore_stage_mem (
    input clk,
    input rst,
    kamacore_pipeline_stage pipeline_ex_mem, 
    kamacore_pipeline_stage pipeline_mem_wb
);
    // Temporarily: Access unmapped SRAM data memory
    // Stage buffer
endmodule
