///////////////
// Writeback //
///////////////

module kamacore_stage_wb (
    kamacore_pipeline_stage pipeline_mem_wb,
    output logic writeback_result
);
    // Decide writeback result
endmodule
