
///////////////////
// Execute stage //
///////////////////

module stage_ex (
    pipeline_stage pipeline_ex
);
    // TODO: Implement 
endmodule