
`import kamacore_pkg::kama_core

///////////////
// Writeback //
///////////////

module stage_wb (
    input logic clk,
    input logic rst,
    kama_core.stage_mem_wb
);
    // TODO: Implement 
endmodule