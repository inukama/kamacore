
module instruction_memory(
);

endmodule