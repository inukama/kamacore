///////////////
// Writeback //
///////////////

module stage_wb (
    pipeline_stage pipeline_wb
);
    // TODO: Implement 
endmodule