
module kama_core(
    input logic clk,
    input logic rst
);



endmodule

