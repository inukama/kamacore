///////////////////////
// Instruction Fetch //
///////////////////////

module kamacore_stage_if (
    input branch_valid,
    kamacore_pipeline_stage pipeline_if_id
);
    // Program counter
    // Access instruction memory
    // Stage buffer
endmodule
