///////////////////
// Execute stage //
///////////////////

module kamacore_stage_ex (
    kamacore_pipeline_stage pipeline_id_ex,
    kamacore_pipeline_stage pipeline_ex_id
);
    // Arithmetic Logic Unit
    // Stage buffer
endmodule
