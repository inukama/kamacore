///////////////////////
// Instruction Fetch //
///////////////////////

module stage_if (
    pipeline_stage pipeline_if
);
    // TODO: Implement 
endmodule