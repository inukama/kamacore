//////////////////
// Memory stage //
//////////////////

module stage_mem (
    pipeline_stage pipeline_mem 
);
    // TODO: Implement 
endmodule