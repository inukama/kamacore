
`import kamacore_pkg::kama_core

///////////////////////
// Instruction Fetch //
///////////////////////

module stage_if (
    input logic clk,
    input logic rst,
    kama_core.stage_if_id
);
    // TODO: Implement 
endmodule