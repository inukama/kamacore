////////////////////////
// Instruction Decode //
////////////////////////

module stage_id (
    pipeline_stage pipeline_id
);
    // TODO: Implement  
endmodule