////////////////////////
// Instruction Decode //
////////////////////////

module kamacore_stage_id (
    input logic clk,
    input logic rst,
    input logic [CPU_WIDTH-1:0] writeback_result,
    kamacore_pipeline_stage pipeline_if_id,
    kamacore_pipeline_stage pipeline_id_ex
);
    // Access register file

    // Generate control signals
    // Stage buffer
endmodule
