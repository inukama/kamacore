
module forwarding_unit();
endmodule
