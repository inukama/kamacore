
`import kamacore_pkg::kama_core

////////////////////////
// Instruction Decode //
////////////////////////

module stage_id (
    input logic clk,
    input logic rst,
    kama_core.stage_if_id,
    kama_core.stage_id_ex
);
    // TODO: Implement  
endmodule