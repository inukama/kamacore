
`import kamacore_pkg::kama_core

//////////////////
// Memory stage //
//////////////////

module stage_mem (
    input logic clk,
    input logic rst,
    kama_core.stage_ex_mem,
    kama_core.stage_mem_wb
);
    // TODO: Implement 
endmodule