
`import kamacore_pkg::kama_core

///////////////////
// Execute stage //
///////////////////

module stage_ex (
    input logic clk,
    input logic rst,
    kama_core.stage_id_ex,
    kama_core.stage_ex_mem
);
    // TODO: Implement 
endmodule