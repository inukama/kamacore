///////////////
// Writeback //
///////////////

module kamacore_stage_wb (
    input clk,
    input rst,
    kamacore_pipeline_stage pipeline_mem_wb,
    output logic [CPU_WIDTH-1:0] writeback_result
);
    // Decide writeback result
endmodule
